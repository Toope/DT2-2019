`include "fir_filter.svh"
bind fir_filter fir_filter_svamod SVA_fir_filter (.*);
bind i2c_slave i2c_slave_svamod SVA_i2c_slave (.*);
