`ifndef SYNTHESIS
timeunit 1ns;
timeprecision 1ps;
`endif

