`include "fir_filter.svh"
///////////////////////////////////////////////////////////////
//
// Template for top-level module
//
///////////////////////////////////////////////////////////////



module fir_filter_svamod
  
  (input logic clk,
   input logic rst_n
   
   );

	
endmodule


